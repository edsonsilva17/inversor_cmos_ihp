** sch_path: /home/edsonihp/ihp130_skel/tarefa1/inversor.sch
.subckt inv vdd out in gnd
*.PININFO out:B vdd:B gnd:B in:B
M1 out in gnd gnd sg13_lv_nmos w=0.45u l=0.15u ng=1 m=1
M2 out in vdd vdd sg13_lv_pmos w=0.9u l=0.15u ng=1 m=1
.ends
.end
